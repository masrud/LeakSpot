b0VIM 7.3      �0T�B� �  masoomeh                                masoomeh-ThinkPad                       ~masoomeh/Research/DevelopedTools/HttpsProxy/node_modules/JSInstrument/lib/JSInstrument.js                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           e                            u       f                     _       �                     d       :                    &       �                    6       �                    m       �             	       W       f             
       ^       �                    P                           ^       k                    X       �                    j       !                    ;       �                    S       �                    \                           	       u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     e       �  p  o     �  �  �  c    �  �  �  �  ]  9    �  �  �  F  E  '        �  �  �  x  c  9  �
  �
  u
  6
  
  �	  �	  �	  K	  	  �  �  �  s  O  I  )  (  �  �  �  �  �  �  ~  b  H      �  d    �  �  �  �  k  X  Q  P  <  ,      �  �  �  �  �  s  O  N  D    �  �  u  Z  >     �  �  �  |  X  W  D    �  �  �                  BlockStatement: 'BlockStatement',         ArrayExpression: 'ArrayExpression',         AssignmentExpression: 'AssignmentExpression',     var Syntax = {      N_LOG_REGEXP_LIT = 44; //RegExp     N_LOG_BUILTIN_DATE = 43,   //Date     N_LOG_BUILTIN_ARRAY = 42,  //Arrays     N_LOG_OBJECT_NEW_INSTANCE = 40, //instances     N_LOG_NULL_LIT = 25,                  N_LOG_UNDEFINED_LIT = 24,     N_LOG_BOOLEAN_LIT = 23,     N_LOG_NUMBER_LIT = 22,     N_LOG_STRING_LIT = 21,        N_LOG_FUNCTION_LIT = 12,  //Function Expression       N_LOG_OBJECT_LIT = 11,   //Object Expression  //anonymous     N_LOG_ARRAY_LIT = 10,   //Array Expression   //anonymous     var        //functions/Builtin Data types.     //Before finalizing and enough testingh let's have the name of the      };         OEXP3: 7         INC: 6,         OEXP2: 5,         PARAMS: 4,         OEXP: 3,         IGNORE: 2,         RHS: 1,     var CONTEXT = {      };         FuncExp: 2         FunctionDec: 1,     var ScopeType = {  //observe function on the specified object.... // If it checks the value of the property, and if it is innerHTML, then it applies //need to handle this during runtime. When a property is being accessed //This is especially true since the name of a property may change. Instead, we  //There is no need for special consideration of innerHTML during instrumentation.      //TODO: take the object that is returned by a function call!     var RP = PREFIX1+"_";     var loggerLib = JSProf;     var PREFIX1 = "JSProf";      //TODO: Callexpression not s      }         this.options.PARSING_MODE = options.parsing_mode;     this.setOptions = function (options) {       // DELETE_INST        : 1,     }         PARSING_MODE       :'PARSE'         LITERAL_INST       : 0,         INFILE_INST        : 0,         RECORD_RIGHT_NULL  : 1, //set to null         ACCUMULATION_POINT : 1, //Reference creation         WRITE_INST         : 1, //Reference creation         ASSIGNMENT_INST    : 1, //Reference creation         MEMBEREXP_INST     : 1,  //ACCESS OBJECT         IDENTIF_INST       : 1,  //ACCESS OBJECT         ARRAYEXP_INST      : 1,  //Create         OBJEXP_INST        : 1,  //Create         PROGRAM_INST       : 1,  //Function Declaration insdie         FUNCDECL_INST      : 1,  //Function Declaration inside         FUNCTINEXP_INST    : 1,  //Create + Function Declaration inside         CALLEXP_INST       : 1,  //ACCESS functions, methods         NEWEXPRESSION_INST : 1,  //Create     this.options = {     //TODO: access to function arguments     var thatModule = this; var JSINSTRUMENT = function(depth) { //module.exports = new (function()   }     return new JSINSTRUMENT(); module.exports = function() {  require('/home/masoomeh/Research/DevelopedTools/HttpsProxy/lib/profilerLib.js'); //var loggerLib = require('../../../lib/profilerLib.js'); var crypto = require('crypto'); var escodegen = require('escodegen'); var esprima = require('esprima'); //var esprima = require('esprima'); var estraverse = require('estraverse'); var fs = require('fs');  //with the default value for this inside a function //inside the logging function, since if it is a this, it will be confused //(a==this), it does not work. Actually, we should not call the object //NOTE:Replacing a[i] = 6 with PE(a,i,6) does not work, since if   //in the code to see what is going wrong!!! //you want to go and dig into the code, then it will be helpful when digging  //In the code, Try to write the beautified version of each file, so that when   // orion.client / bundles / org.eclipse.orion.client.javascript / web / javascript / contentAssist / esprimaVisitor.js  //general AST traversal ad    Q     	       �  �  �  �  c  U  S  R  Q  P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     }             }                 return newCode;                 var newCode = escodegen.generate(ast, codegenerateoptions );                       }, parse: esprima.parse}; ad  #        u       �  �  ~  Z  "  �  �  �  j  6    �  �  �  ^  :    �  �  �  j  <       �  �  x  V  ,    �
  �
  �
  N
  
  �	  �	  �	  �	  �	  u	  o	  n	  H	  	  	  	  �  �  �  �  �  �    g  L  2  	  �  �  �  �  �  �  �  n  .  '  &    �  �  �  �    d  A  7    �  �  �  �  �  {  U  G  =  )  #    �  �  �    @  ?    �  �  �  �  �  �  W    �  �  �  �  �  d  Z  M  1  0                                                 ret = replaceInExpr(              lid = getLId();         else         }             lid = getPreviousLId();         if (ReUseLId) {             logFunction = logFuncName;         if (logFuncName !== undefined)         var ret;         var lid;         var logFunction= logFunctionName ( loggerLib.consts.logRead );     function wrapRead(node, logFuncName, ReUseLId) {      }         return ret;         );         body             "\n try{"+RP+"1}\n catch (e) \n{ }\n finally \n{ JSProf.FLUSH(); }\n",         var ret = replaceInStatement(n_code+          var n_code = '\n    require("'+preFile+'");\n' + '\n';          var preFile = path.resolve(__dirname,'../../../lib/profilerLib.js');         var path = require('path');     function prependScriptBody(node, body) {          }         return res;         }             }                 res[i] = fun(arr[i]);             if (i in arr) {         for (var i = 0; i < len; i++) {         var res = new Array(len);          }             throw new TypeError();         if (typeof fun != "function") {         }             throw new TypeError();         if (!isArr(arr)) {         var len = arr.length;     function MAP(arr, fun) {      }         return Object.prototype.toString.call( val ) === '[object Array]';     function isArr(val) {      };         return Object.prototype.hasOwnProperty.call(obj, prop);     function HOP(obj, prop) {      }         return createLiteralAst(tempIid);         var tempIid = LID - inc;     function getPreviousLId() {      }             return createLiteralAst(tmpIid);         LID = LID + inc;          var tmpIid = LID;      function getLId() {      var LID = 1+inc;     var inc = 1;       }         return {type: Syntax.Identifier, name: name};     function createIdentifierAst(name) {      }         return {type: Syntax.Literal, value: name};     function createLiteralAst(name) {      }         return PREFIX1+"."+funcname;     function logFunctionName(funcname) {      };         WithStatement: 'WithStatement'         WhileStatement: 'WhileStatement',         VariableDeclarator: 'VariableDeclarator',         VariableDeclaration: 'VariableDeclaration',         UpdateExpression: 'UpdateExpression',         UnaryExpression: 'UnaryExpression',         TryStatement: 'TryStatement',         ThrowStatement: 'ThrowStatement',         ThisExpression: 'ThisExpression',         SwitchCase: 'SwitchCase',         SwitchStatement: 'SwitchStatement',         SequenceExpression: 'SequenceExpression',         ReturnStatement: 'ReturnStatement',         Property: 'Property',         Program: 'Program',         ObjectExpression: 'ObjectExpression',         NewExpression: 'NewExpression',         MemberExpression: 'MemberExpression',         LogicalExpression: 'LogicalExpression',         LabeledStatement: 'LabeledStatement',         Literal: 'Literal',         IfStatement: 'IfStatement',         Identifier: 'Identifier',         FunctionExpression: 'FunctionExpression',         FunctionDeclaration: 'FunctionDeclaration',         ForInStatement: 'ForInStatement',         ForStatement: 'ForStatement',         ExpressionStatement: 'ExpressionStatement',         EmptyStatement: 'EmptyStatement',         DebuggerStatement: 'DebuggerStatement',         DoWhileStatement: 'DoWhileStatement',         ContinueStatement: 'ContinueStatement',         ConditionalExpression: 'ConditionalExpression',         CatchClause: 'CatchClause',         CallExpression: 'CallExpression',         BreakStatement: 'BreakStatement',         BinaryExpression: 'BinaryExpression', ad  J   �     _       �  �  �  �  �  �  �  X  7  �  �  c  R  G  3  -  ,  �  �  �  �  �  p  `  U  A  ;  :    �    m  ?  .  #    	    �  �  j  3      �
  �
  �
  �
  �
  �
  t
  F
  
  �	  �	  �	  �	  �	  '	  �  �  �  e    �  �  �  �  _  ^    �  U  �  �  K  J  I  $  �  �  k  J  +    �  �  �  �  �  I  �  �  <  �  �                                                                                            else if (actionType === logFunctionName( loggerLib.consts.logPutDotNull))                     actionType = logFunctionName( loggerLib.consts.logPutFieldBracket );                 else if (actionType === logFunctionName( loggerLib.consts.logPutFieldDot) )                     actionType = logFunctionName( loggerLib.consts.logGetFieldBracket);                 if (actionType == logFunctionName( loggerLib.consts.logGetFieldDot))             else {             }                 return ret;                  );                     node.property                     node,                     nproperty,                     node.object,                     getLId(),                     //actionType+"("+RP+"1, "+RP+ "2, "+RP+"3)["+RP+"4]",                     actionType+"("+RP+"1, "+RP+ "2, "+RP+"3, "+RP+"4)["+RP+"5]",                 ret = replaceInExpr(                       actionType = logFunctionName( loggerLib.consts.logPutBracketNull);                 else if (actionType === logFunctionName( loggerLib.consts.logPutDotNull))                     actionType = logFunctionName( loggerLib.consts.logPutFieldBracket );                 else if (actionType === logFunctionName( loggerLib.consts.logPutFieldDot))                     actionType = logFunctionName( loggerLib.consts.logGetFieldBracket);                 if (actionType == logFunctionName( loggerLib.consts.logGetFieldDot ))                      nproperty = createLiteralAst(node.property.name);                 else                 }                     }                         //console.log("************");                         nproperty = createLiteralAst(node.property.value);                      if (node.property.type == 'Literal') {                 if ( node.property.name == undefined) {                 var nproperty;                 //return node; //TODO: FIX THIS             if ( ( node.property.type === "Identifier" ) || ( node.property.type === 'Literal' ) ) {         if ( node.computed == true) {     function wrapGetPutField(node, actionType) {      }         return sha1.digest("hex").toString("utf8");         sha1.update(new Buffer(tname));         var sha1 = crypto.createHash("sha1");         var tname = node.object.type + "-" + node.object.name;     function makeTempVar(node) {      }         return ret;         );             node             tret,             getLId(),             logFuncName+"("+RP+"1, "+RP+"2, "+RP+"3)",         var ret = replaceInExpr(         var tret = wrapIW(createIdentifierAst(lhs.name));     function wrapWriteWithUndefinedCheck(node, lhs, logFuncName) {      }         return ret;         );             node             createIdentifierAst("undefined"),             node,             logFunctionName ( loggerLib.consts.logUndefined ) + "(typeof " +  RP+"1" + " === 'undefined' ?"+RP+"2: "+RP+"3)",         var ret = replaceInExpr(     function wrapIW(node) {      }         return ret;         );             val             lhs,             getLId(),             logFuncName+"("+RP+"1, "+RP+"2, "+RP+"3)",         ret = replaceInExpr(         var ret;     function wrapWrite(val, lhs, logFuncName) {      }         return ret;         );             node             createIdentifierAst("undefined"),             getLId(),             logFunctionName( loggerLib.consts.logReadUndefined ) + "("+ RP+ "1, typeof " +  node.name + " === 'undefined' ?"+RP+"2: "+RP+"3) ",         var ret = replaceInExpr(     function wrapReadWithUndefinedCheck(node) {      }         return ret;         );             node              lid,             logFunction+"("+RP+"1, " +RP+"2)", ad  %   �     d       �  �  t  9    �  �  �    V  �  �  �  t  L  !  �  �  �  �  �  �  g  $  
  �  �  �  �  r  Y  O  I  H  $    �
  �
  �
  ?
  
  
  �	  �	  �	  Q	  	  �  �  �  �         �  �  �  v  >  !      �  n  R  H  9           �  �  �  1    �  �  A    �  �  �  �  �  �  �  K  :    �  �  �  w  c  ]  Z  )    �  �                                               if (scope.hasVar(node.left.name)) { // if a is already defined         var ret;     function instrumentIdentifierSetNull(node) {        }         return ret;         }                ret = wrapRead(node.right,logFunctionName( loggerLib.consts.logGlobalVar));         } else {              ret = node.right;          if (scope.hasVar(node.left.name)) {          var ret;     function instrumentGlobalVariableReference(node) {          }         //return ret;         //}         //    return node;         //} else {         //    var ret = instrumentLoad(node.left);         //if (node.left.type === 'Identifier') {         //to apply instrumentLoad function with a different parameter.         //difference is that the object is also being read. I just need         // It can be treated as a write, since it is written. The only          //at the moment.         //we are not targetting number objects, so we skip wrting this function         //Actually since all of the other operators are used on number, and          return node;     function instrumentLoadModStore(node) {      }         }             return node;         else {         }                 return ret;                 ret = wrapGetPutField(node, logFunctionName( loggerLib.consts.logGetFieldDot));         else if ( node.type === 'MemberExpression' ) {         }             }                     return ret;                  ret = wrapReadWithUndefinedCheck(node);             } else {                 return ret;                  ret = wrapRead(node);             } else if (scope.hasVar(node.name)) {                 return node;              node.name === "eval" || node.name === "arguments"){ //Last Condition is for Facebook             } if(node.name === PREFIX1 ||                     return node;                 else                 }                     return ret;                      ret = wrapLiteral(node, N_LOG_NUMBER_LIT);                 if (thatModule.options.LITERAL_INST==1) {              } else if (node.name === "NaN" || node.name === "Infinity") {                     return node;                 else                 }                     return ret;                      ret = wrapLiteral(node, N_LOG_UNDEFINED_LIT);                 if (thatModule.options.LITERAL_INST==1) {              if (node.name === "undefined") {         if (node.type === 'Identifier') {         var ret;     function instrumentLoad(node) {      }         }             return ret;              );                 node.property                 //node,                 createLiteralAst(node.property.name),                 node.object,                 getLId(),                 actionType+"("+RP+"1, "+ RP+"2, "+RP+"3)."+RP+"4",             ret =  replaceInExpr(         else {         }             }                     return ret;                      );                         createIdentifierAst (hashedname)                         tret.arguments[0],                         node.property,                          createIdentifierAst (hashedname),                         node.object,                         getLId(),                         actionType+"("+RP+"1, "+RP+ "2, "+RP+"3 = "+RP+"4, "+RP+"5) ["+RP +"6]",                     ret = replaceInExpr(                      createIdentifierAst (hashedname));                     node.object,                     actionType+"("+RP+"1[ "+RP+ "2])",                 var tret = replaceInExpr(                 hashedname = PREFIX1+".TMPS.t"+hashedname;                 var hashedname = makeTempVar(node);                      actionType = logFunctionName( loggerLib.consts.logPutBracketNull); ad  A	  �	     &       �  �  x  2  �  �  �  �  �  �  v  /  �  �  v  3  �  �  �  �  E  �  �  �  �  �  �  �  a  �
  �
  ~
  j
  d
  c
  >
  ,
  �	  �	  �	  p	  L	  8	  	  �  �  �  O  ,    
  	  �  z  :      �  �  �  �  x  *  	  �  �  �  L  �  �  �  �  f  E  �  �  �  �  \    �  r  T    �  �  �  �  �  �  �  �          function getPropertyAsAst(ast) {       }         }                 return node;              }                 node.right = ret;                 ret = instrumentAccumulationPoint(node, ReUseLId);                 // right one.                 // left side and the object on the right side by wrapping the                  // TODO in script to process data: connect the container on the                 // get the iid of the left side and use that for the right             if ( (thatModule.options.ACCUMULATION_POINT==1) && (rightType===true)) {              }                 node.left = ret;                 ret = wrapGetPutField(node.left, logFunctionName(loggerLib.consts.logPutFieldDot));                 ReUseLId = true;             else if (thatModule.options.WRITE_INST===1) {             }                 }                     node.left = ret;                     ret = wrapGetPutField(node.left, logFunctionName(loggerLib.consts.logPutDotNull));                 if (thatModule.options.RECORD_RIGHT_NULL===1) {                 rightType = false;             if ((node.right.type==="Literal")&&(node.right.value===null))  {                          // it is set to Null             //TODO: remove the following, later add support for the case that             var rightType=true;             var ReUseLId = false;         } else {  //a.b =              return node;                  }                  }                     node.right = ret;                     ret = instrumentIdentifierSetNull(node);                     if ((node.right.type==="Literal")&&(node.right.value===null))  {              if (thatModule.options.RECORD_RIGHT_NULL===1) {               }                  }                  node.right = ret;                  ret = instrumentWriteToIdentifier(node);                 else {                 }                 if ((node.right.type==="Literal")&&(node.right.value===null)) {              if (thatModule.options.WRITE_INST===1) {             // }                //    node.right = ret;             //    ret = instrumentGlobalVariableReference(node);             //if (thatModule.options.GLOBAL_VAR        return node;         if (node.left.type === 'Identifier') { // a =          var ret;      function instrumentStore(node) {      }         return ret;             ret = wrapRead(node.right, logFunctionName( loggerLib.consts.logRightSidePutDot), ReUseLId);         else             ret = wrapRead(node.right, logFunctionName( loggerLib.consts.logRightSidePutBracket), ReUseLId);         if (node.left.computed==true)         var ret;     function instrumentAccumulationPoint(node, ReUseLId) {      }         return ret;         }                    logFunctionName( loggerLib.consts.logWriteUndefined));                ret = wrapWriteWithUndefinedCheck(node.right, node.left,              //THIS WOULD MEAN A GLOBAL REFERENCE              //it is inside a variable declaration             //generated code. Note that ' var a = ..' is OK. since              //and if it is not defined results in an error in the          } else { // if a is not defined. Since JSRecord.Write calls a                  logFunctionName( loggerLib.consts.logWrite));             ret = wrapWrite(node.right, node.left,          if (scope.hasVar(node.left.name)) { // if a is already defined         var ret;     function instrumentWriteToIdentifier(node) {          }         return ret;         }                    logFunctionName( loggerLib.consts.logWriteUndefinedNull));                ret = wrapWriteWithUndefinedCheck(node.right, node.left,          } else {                  logFunctionName( loggerLib.consts.logWriteNull));             ret = wrapWrite(node.right, node.left,  ad     �     m       �  �  �  �  -    �  �  g  <  	  �  �  �  e  S  D  C    �  y  <  &    �  �  �  �  �  c  G  A  @    �
  �
  �
  �
  r
  
  �	  �	  ^	  D	  .	  	  �  �  �  �  �  U  F     �  �  �  N  0       �  �  �  �  �  >  (      �  �  �  �  �  �  O      	  �  �  �  U  #  �  �  �  |  r  h  O  E  D  �  �  �  �  �  n  U  S  =  7  6  5  �  �  �  �                  // arguments, length, keys     //TODO, do the same for access to native properties!        }         return false;               return true;         if (node.callee.name === "setTimeout")   //for Facebook          }             return true;         {         if ( (node.callee.type==='MemberExpression') && ( (node.callee.property.name === 'bind')  )   )          }             return true;         {         )         )         (node.callee.property.name === 'require')          (node.callee.property.name === 'inherits') ||         ( (node.callee.property.name === 'base')||          (node.callee.object.name === 'goog') &&           if ( (node.callee.type==='MemberExpression') &&         }*/             //ret = wrapNewExpression(node, 'objcreate'); //TODO: wrap object.create()             return true;         {          )         (node.callee.property.name === 'create')         (node.callee.object.name === 'object') &&         /*if ( (node.callee.type==='MemberExpression') &&      function stopInstrumentingCallExpression(node) {       }         return ret;         );             ast             getLId(),             logFunctionName( loggerLib.consts.logFuncCall) +"("+RP+"1, "+RP+"2, "+(isCtor?"true":"false")+")",         var ret = replaceInExpr(     function wrapFunCall(ast, isCtor) {      }         }             return ret;              );                  node.property                 createLiteralAst(node.property.name),                 base,                 getLId(),                 logFunctionName( loggerLib.consts.logMethodCall) + "("+RP+"1,  "+RP+"2, "+RP+"3)."+RP+"4",              var ret = replaceInExpr(          else {         //TODO: handle the case where node.computed === false, e.g., a[i++]()         }             return ret;              );                 property                 createLiteralAst(type),                 offset,                 base,                 getLId(),                 logFunctionName( loggerLib.consts.logMethodCall) + "("+RP+"1, "+RP+"2, "+RP+"3, "+RP+"4)["+RP+"5]",              var ret = replaceInExpr(              var type=1;         if (node.computed === true ) { //TO handle cases such as a[0]() which happened in google     function wrapMethodCall(node, base, offset , property, isCtor) {      }         return ret[0].expression;         var ret =  replaceInStatement.apply(this,arguments);     function replaceInExpr(code) {      }         return newAst.body;         var newAst = transformAst(ast, visitorReplaceInExpr, undefined, undefined);         var ast = esprima.parse(code);          }             }                 return node;                 }                     }                         node.body = node.body[0].expression;                     if (node.body[0].type === 'ExpressionStatement' && isArr(node.body[0].expression)) {                 if (node.body[0] != undefined) {             'BlockStatement' : function(node) {              },                 }                     return node;                 } else {                     return asts[i];                     var i = parseInt(node.name.substring(RP.length));                 if (node.name.indexOf(RP) === 0) {             'Identifier': function(node) {         var visitorReplaceInExpr = {         //its value later when it is being called         //Here asts in a closure, that's why the visitorReplaceInExpr can access         var asts = arguments;         //Here is the part for making the part that is needed to be added to the AST.     function replaceInStatement(code) {      }         return ast.computed?ast.property:createLiteralAst(ast.property.name); ad     �     W       �  r  q  $  �  �  a  `    �  �  �  }  =  �  �  �  �  6  �  �  �  N    �
  �
  q
  6
  (
  '
  �	  �	  i	  	  �  j  G      �  �  i  %  �  �  �  �  r  q  p  B  A  �  �  �  �    �  �  �  �  Y  G  A  @      �  �  �  r  $  �  �  �  �  �  p  _  3        
  �  �  �  �                                       var ret = replaceInExpr( RP+"1 "+op+" "+RP+"2",          function wrapRHSOfModStore(node, left, right, op) {      }         }             return ret;             ret = wrapFunCall(ast, isCtor);         } else {             return ast;         } else if (ast.type ==='Identifier' && ast.name === "eval") {              }                 return ret;                     ast.property, isCtor);                 ret = wrapMethodCall(ast, ast.object, getPropertyAsAst(ast),              else {                 return ast;             if (checkToInstrument(ast,0) == 1) //TODO         if (ast.type==='MemberExpression') {         var ret;     function instrumentCall(ast, isCtor) {      }         return 0;         //console.log(node.property.name);         }             return 1;         ){         ( (node.object.name==="window") && (node.property.name==="postMessage") )         ( (node.object.name==="Math") && ( (node.property.name==="random")|| (node.property.name==="floor") || (node.property.name==="pow"))) ||         if ( ( (node.object.name==="console") && (node.property.name==="log") ) ||              return 1;         if (NoInstrumentNoChange.indexOf( node.property.name ) >=0 )      function checkToInstrument(node, level) {       // 'toString', 'removeChild', 'pop'     // 'appendChild',     // 'getElementById', 'createElement',     ];         'isDisposed', 'toString', '_DumpException', 'dispatchEvent'         'concat', 'toLowerCase', 'split', 'unshift', 'toUpperCase',         'insertBefore', 'charAt', 'substring', 'clearTimeout',     var NoInstrumentNoChange=['toLocaleString', 'exec', 'getElementsByTagName',     //TODO: make this list complete      //This is even true for push and get.     //perform the instrumentation.     // It is using the definition by the program. although this means that we need to      // this means that this function is defined by the program, otherwise, it means that     // If when referencing to this function, the object id is created before,      // isCollapsed, dispatchEvent in Gmail.     // creates a new Definition. For example, I have seend for the      // For some functions, event though it is a native function, the program       'apply'];         'create', 'caller', 'constructor', 'call', 'bind',         'freeze', 'defineProperty', 'defineProperties',          'getOwnPropertyNames', 'getOwnPropertyDescriptor',         'hasOwnProperty', 'is', 'getPrototypeOf',          'isPrototypeOf', 'isFrozen', 'isExtensible',          'preventExtensions', 'name', 'isSealed',          'prototype', 'propertyIsEnumerable',          'toString', 'toLocaleString', 'seal', 'getSelection', 'isCollapsed',          'setRequestHeader', 'setTimeout', 'clearTimeout',         'addEventListener', 'attachEvent', 'preventDefault', 'send', 'error', 'match','open',         'dispatchEvent', 'toLowerCase', 'focus',         'slice',  //Array         'charAt',         'queryCommandSupported', 'getElementsByTagName',              //DOM         'createTextNode', 'createElement', 'execCommand', //DOM         'getTime', //Date         'exec',   //RegExp         'indexOf', 'unshift',         'get', 'join', 'split', 'getElementById', 'valueOf',      var NoInstrumentPropertiesName=['replace', 'call', 'apply', 'substr', 'push',      //is much higher than size overhead.     //Actually in the profilerLib is more important. Since the network overhead     //those issue that mentioned in that ECOOP paper about object.create!     //TODO: add this point to the paper that by dynamic analysis, we resolve      //sent to the proxy. This reduces the communication overhead.     //TODO: Also do this during runtime, so that the info for these are not ad  J   �     ^       �  �  �  �  x  I  %  �  �  �  |  m  U  K  B    �  �  l  W  )      �  �  �  �  @  &    �  �  �  �  �  �  �  [  �
  �
  b
  a
  H
  >
  =
  
  
  �	  k	  Q	  <	  '	  	  	  �  �  �  �  �  �  >  =    �  �  �  q  b  a  I  ?  >  �  �  �  b  E    �  �  b  &  �  �  g    �  �  1  �  �  �  2  �  �                                                                                                                                estraverse.traverse(thisnode, {                                                     console.log('...........');                                                      var testUsedinFunc=false;                                                 if (scope.vars[thisnode.id.name] === "defun") {                                             if (scope.vars[thisnode.id.name] !== undefined) {                                             console.log(scope.vars);                                             console.log(thisnode.id.name);                                             console.log(thisnode.type);                                         {                                         if ((thisnode.type == 'FunctionDeclaration'))                                     enter: function(thisnode){                                 estraverse.traverse(node, {                                 console.log("name...."+name);                             if (scope.vars[name] ==="var") {                         if (HOP(scope.vars, name)) {                     for (var name in scope.vars) {                 if (scope) {                 //TODO: complete implenting context refences             var ret = [];         function syncCreateRef (node, scope, isScript) {     //TODO: closure reference should be done on function arguments as well.          }             return ret;              );                 val                 //name,                 getLId(),                 logFunctionName( loggerLib.consts.logFuncDeclaration)+"("+RP+"1, "+RP+"2 )",             var ret =replaceInStatement(              //name is added in the above to differentiate betweeen functions allocated within a scope         function createCallInitAsStatement(node, name, val, isArgumentSync) {            }             return ret;              );                 func                 val,                 getLId(),                 logFunctionName( loggerLib.consts.logCreateContextReference )+"("+RP+"1, "+RP+"2, "+RP+"3)",             var ret =replaceInStatement(          function createContextReference(node, val, func) {          }             return ret2;              node.argument, ret);             var ret2 =  replaceInExpr( RP+"1 =  " + logFunctionName( loggerLib.consts.logWrite)  +"( "+RP+"2 )",             var ret = wrapRHSOfModStore(node, node.argument, right, node.operator.substring(0,1)+"=");             var right = createLiteralAst(1);         function instrumentPreIncDec(node) {          }             return ret;              );                 createLiteralAst(funId)                 node,                 getLId(),                 logFunctionName( loggerLib.consts.logLiteral)+"("+RP+"1, "+RP+"2, "+RP+"3)",             var ret =  replaceInExpr(         function wrapLiteral(node, funId) {                  }             return ret;             );                 createLiteralAst(objTypeName)                 ast,                 getLId(),                 logFunctionName( loggerLib.consts.logNewObject)+"("+RP+"1, "+RP+"2, "+RP+"3)",             var ret =  replaceInExpr(         function wrapNewExpression(ast, objTypeName) {                  }             return ret;             );                 ast                 getLId(),                 logFunctionName( loggerLib.consts.logCallExp) +"("+RP+"1, "+RP+"2)",             var ret =  replaceInExpr(         function wrapCallExp(ast) {         //case of renaming this does not hold.         //TODO: Identify the name of function that is wrapped, although in          }             return ret;             left, right); ad     w     P       �  5  �  �  �  m  l  $  �  g    �  �  k  A  �  �  �  q  S  R    �
  m
  (
  '
  �	  �	  [	  	  	  �  �  \  �  �  �  a    �  �  �  j  i  3  �  �  l  J  I  $    �  �  �  �  �  �  �  �  |  _  S  R      �  �  t  B  *      �  �  �  R    �  w  v                                                             ret = ret.concat(createCallInitAsStatement(node,                                 //ident.loc = scope.funLocs[name];                                 var ident = createIdentifierAst(name);                             if (scope.vars[name] ==="defun") {                         if (HOP(scope.vars, name)) {                     for (var name in scope.vars) {                 if (scope){                  }*/                 true));                 createIdentifierAst("arguments"),                 createLiteralAst("arguments"),                 ret = ret.concat(createCallInitAsStatement(node,             /* if(!isScript) {             var ret = [];         function syncDefuns(node, scope, isScript) {          }                   return ret;                  }                      }                         }                            } */                                  }                                 }                                 }                                     }                                 createIdentifierAst(name)));                                 //createLiteralAst(name)));                                 ret = ret.concat(createContextReference(node,                                 if (testUsedinFunc) {                                  });                                 }                                 }                                 createIdentifierAst(name))); //*                                 ret = ret.concat(createContextReference(node,                                 /* console.log("***************");                                 testUsedinFunc=true;                                 {                                 if ((thisnode.type == 'Identifier')&& (thisnode.name===varname))                                 enter: function(thisnode){                                 estraverse.traverse(node, {                                 var testUsedinFunc=false;                                  if ( parentScope.vars[varname] === "var" ) {                                 for (var varname in parentScope.vars) {                                 if (parentScope!==null) {                                 var parentScope = scope.getParentScope();                                  //and applycontex reference to them.                                 //get the local variables of the parent scope                                 //check to see if the function closes over any variable                             /*if (scope.vars[name] ==="var") {                              }                                 });                                     }                                         }                                         else if ((thisnode.type == 'FunctionExpression')) {                                         }                                             }                                                 }                                                         ));                                                              createLiteralAst(thisnode.id.name)                                                             createIdentifierAst(name),                                                         ret = ret.concat(createContextReference(node,                                                     if (testUsedinFunc)                                                      });                                                         }                                                                  testUsedinFunc=true;                                                             if ((thenode.type == 'Identifier')&& (thenode.name===name))                                                         enter: function(thenode) { ad  >   �     ^       �  T  )     �  �  �  �  �  P    �  �  �  b    �  �  �  d  F  ,    �  �  �  �  �  �  �  �  �  l  K    �
  �
  �
  �
  �
  �
  ^
  =
  (
  
  �	  �	  �	  `	  $	  �  �  �  o  8  �  �  �  [  4    �  �  �  J  &  	  �  �  �  �  �  �  �  h  .  �  �  �  v  '  �  �  g  )    �  �  �  �  �  h     �  �                                                                                // What about accesses. Here a write happend, but we are not                  // TODO: any reference is created here? global, local?              'VariableDeclaration': function (node) {                },                 return node;                 scope = scope.parent;                 }                     node.body = ret;                     ret = prependScriptBody(node, node.body);                     //instrumented file                     //content of profilerLib.js to the beginnign of the                      //commented. To run in local mode, we need them to add the                     //To run in Proxy mode, the following two lines should be                  if (thatModule.options.INFILE_INST == 1) {                 }                     node.body = ret;                     ret = instrumentScriptEntryExit(node, node.body);                 if (thatModule.options.PROGRAM_INST==1) {                 var ret;              'Program': function(node) {              },                   }                     }                         return node;                     } else {                         return ret;                         var ret = wrapLiteral(node, litType);                         }                                   break;                                 litType = N_LOG_BOOLEAN_LIT;                             case 'boolean':                                 break;                                     litType = N_LOG_REGEXP_LIT;                                 else                                      litType = N_LOG_NULL_LIT;                                 if (node.value === null)                             case 'object': // for null                                 break;                                 litType = N_LOG_STRING_LIT;                             case 'string':                                 break;                                 litType = N_LOG_NUMBER_LIT;                             case 'number':                         switch(typeof node.value) {                         var litType;                     if (context === CONTEXT.RHS){                 {                 else                     return node;                 if (thatModule.options.LITERAL_INST == 0)              'Literal': function(node, context) {         var visitorRRPost = {          }             'FunctionExpression': setScope             'FunctionDeclaration': setScope,             'Program': setScope,         var visitorRRPre = {          }             scope = node.scope;         function setScope(node) {          var scope;          }                     return ret;                  }                         }                             }                                 } */                             false));                             createIdentifierAst(name),                             createLiteralAst(name),                             ret = ret.concat(createCallInitAsStatement(node,                             if (scope.vars[name] ==="var") {                             }                                 true));                             createIdentifierAst(name),                             createLiteralAst(name),                             ret = ret.concat(createCallInitAsStatement(node,                         /*       if (scope.vars[name] ==="arg") {                               }                                  false));                                     ident,                                     //wrapLiteral(ident, ident, N_LOG_FUNCTION_LIT), //No Need to wrap this one                                     createLiteralAst(name), ad     �     X       �  e    �  t  +  �  �  i    �  �  �  �  y  \  M  L    �  �  �  �  E    �
  �
  s
  ?
  >
  �	  �	  �	  �	  v	  u	  t	  E	  ,	  �  �  �  {  4      �  �  q  L  �  �  �  �  �  �  �  P    �  �  �  �  X  B  )  �  �  �  �  q  >    �  �  �  �  5  �  �  �  �    K    �  �  �  �                                    }                     return node;                     scope = scope.parent; //TODO: what's the use of this!!!!!!                 if (thatModule.options.FUNCDECL_INST==0) {             "FunctionDeclaration": function(node) {             },                 }                     return ret;                     scope = scope.parent;                     var ret = wrapNewExpression(node, N_LOG_FUNCTION_LIT);                     node.body.body = instrumentFunctionEntryExit(node, node.body.body);                 else {                 }                     return node;                     scope = scope.parent;                 if (thatModule.options.FUNCTINEXP_INST==0) {             'FunctionExpression': function(node) {             //TODO: monitor function arguments as accesses             },                 }                     return ret;                         ret = instrumentLoadModStore(node);                     else                     }                         ret = instrumentStore(node);                     if ( node.operator === "=" ) {                     var ret;                 else {                     return node;                 if (thatModule.options.ASSIGNMENT_INST==0)             'AssignmentExpression': function(node) {              },                 return ret;                 }                     ret = node;                     }                         node.arguments = MAP(node.arguments, wrapEvalArg); // TODO                         return node;                     if (isEval) {                     node.callee = callee;                     var callee = instrumentCall(node.callee, false);                      node.callee.name === "eval";                     var isEval = node.callee.type === 'Identifier' &&                  else {                 }                         ret = node;                if ((thatModule.options.CALLEXP_INST==0)||(stopInstrumentingCallExpression(node))) {                 var ret;             "CallExpression": function(node) {               },                 }                     return ret1;                     var ret1 = wrapNewExpression(node, objKind);                     node.callee = instrumentCall(node.callee, true);                          objKind = node.callee.type;                     else                          objKind = N_LOG_OBJECT_NEW_INSTANCE                     else if (node.callee.type == 'MemberExpression')                             objKind = node.callee.name                     if ( node.callee.type == 'Identifier' )                     var objKind;                 else {                         return node;                 if (thatModule.options.NEWEXPRESSION_INST == 0)             'NewExpression': function(node) {              },                 return node;                 node.declarations = declarations;                 });                     return def;                     }                         def.init = init;                         var init = def.init; //TODO: call wrapWrite here.                      if (def.init !== null) {                 var declarations = MAP(node.declarations, function(def){                 // an assignment expression without a variable declaration.                 // so, we need to add references that are created using                  // is considered a global reference. Please note that in doing                  //into scope variable. If the parent of a scope is null then it                 // knowing whether it is a global reference or not needs looking                 // if it is a global reference, then  it adds a reference.                  // monitoring writes. local references are not monitored. Only ad     �     j       �  �  g  E  3  $  �  �  �  �  6      �  �  �  �  i  0    �  �  �  x  i  h  4  �  �  �  �  U  0    �
  �
  �
  �
  �
  �
  V
  
  �	  �	  �	  u	  Q	  4	  	  �  �  �  �  �  �  O  +    �  �  �  �  b  E  7  -  ,  �  �  �  �  �  Q    �  �  �  �  n  U  K  J      �  k  C    �  �  �  �  W  )  �  �  �  �  `  =  +  
  �  �  �  �  �                                }             return ret;             }                 else return ret;                 }                     return ret[0];                     //console.log(ret[0]);                     );                         node.left                         getLId(),                         logInnerHTMLObserver+"("+RP+"1, "+RP+"2)",                     ret = replaceInStatement(                 if (node.left.property.name === "innerHTML") {                                   console.log("...................");                 console.log(node.left.property.name);                 console.log(node.left.property);                 console.log(node.left);                 //test to see if the property name can be changed TODO             if ((node.type === "AssignmentExpression")&&(node.operator==="=")) {             var ret=[];         /*function createNewStatement(node ) {          }             return body;             //body = t3.concat(ast);             //var t3 = syncCreateRef(node, scope, false);             //TODO: update this later:              var body = t2.concat(ast);             var t2 = syncDefuns(node, scope, false);         function   instrumentFunctionEntryExit (node, ast) {          }             return ret;             var ret = syncDefuns(node, scope, true).concat(body);         function instrumentScriptEntryExit(node, body) {          }             }                 return node;                 //node.argument = ret;                 //var ret = instrumentLoad(node.argument);            'ReturnStatement': function(node) {                         },                 return node;                 //node.right = ret;                 //var ret = instrumentLoad(node.right);                 //TODO            'ForInStatement': function(node) {                         },                 }                     }                         return node;                     } else {                         return ret;                         var ret = instrumentLoad(node);                     if (context === CONTEXT.RHS) {                 else {                         return node;                 if (thatModule.options.MEMBEREXP_INST==0)            'MemberExpression': function(node, context) {                         },                    }                     }                             return node;                     else {                     }                          return ret;                          var ret = instrumentLoad(node);                     if (context === CONTEXT.RHS){                 else {                         return node;                 if (thatModule.options.IDENTIF_INST==0)              'Identifier': function(node, context) {              },                 }                     return ret1;                     var ret1 = wrapNewExpression(node, N_LOG_ARRAY_LIT);                 else {                         return node;                 if (thatModule.options.ARRAYEXP_INST==0)             "ArrayExpression": function(node) {             },                 return node;             "UnaryExpression":function(node) {             },                 }                     return ret1;                     var ret1 = wrapNewExpression(node, N_LOG_OBJECT_LIT);                 else {                         return node;                 if (thatModule.options.OBJEXP_INST==0)             "ObjectExpression": function(node) {             },                 }                     return node;                      scope = scope.parent;                     node.body.body = instrumentFunctionEntryExit(node, node.body.body);                 else { ad  |   �     ;       �  �  �  J    �  �  7    �  �  �  �  �  ~  f  Z  Y    �  �  �  �  x  C  B    �  ~  T  )  �
  �
  0
  �	  t	  ?	  �  c  �  �  8  �    �  5  �  d    �  a    �  a    �  �  �  �  �                                                                                                                                                              }                                     newContext = CONTEXT.IGNORE;                                  ) {                                     || (type === 'BreakStatement' && key ==='label')                                     || (type === 'ContinueStatement' && key ==='label')                                     || (type === 'LabeledStatement' && key ==='label')                                     || (type === 'CatchClause' && key ==='body')                                     || (type === 'CatchClause' && key ==='param')                                     || (type === 'NewExpression' && key === 'callee'  )                                     || (type == 'ThrowStatement' && key === 'argument' )                                     || (type === 'UnaryExpression' && key === 'argument' && node.operator === 'delete')                                      || (type === 'VariableDeclarator' && key === 'id')                                      || (type === 'MemberExpression' && node.computed && key === 'property')                                     || (type === 'MemberExpression' && node.computed && key === 'object')                                     || (type === 'MemberExpression' && !node.computed && key === 'object') //TODO: why did you add these two lines at first!!! It is related to wrapGetPutField                                     || (type === 'MemberExpression' && !node.computed && key === 'property')                                     || (type === 'ForInStatement' && key === 'left')                                      || ((type === 'FunctionDeclaration') && key === 'id')                                     || ((type === 'FunctionExpression' || type === 'FunctionDeclaration') && key === 'id')                                     (node.callee.type === 'Identifier' && node.callee.name === 'eval')))                                 (node.callee.type === 'MemberExpression' || node.callee.type === 'Identifier'  ||                                  key === 'callee' &&                                  || ( (type === 'CallExpression' || type === 'NewExpression') &&                                      || (type === 'UpdateExpression' && key === 'argument')                                 if ( (type === 'AssignmentExpression' && key === 'left')                              //if ( type === 'MemberExpression' && node.computed )                         if (typeof child === 'object' && child !== null ) {                          child = node[key];                                 continue;                             if (type === 'Property' && ( node.kind === 'get' || node.kind=== 'set' ) )                     if (node.hasOwnProperty(key)) {                  for (var key in node) {                      visitorPre[type](node, context);                 if (visitorPre && HOP(visitorPre,type))                   type = node.type;                   var key, child, type, ret, newContext;             function transformAst(node, visitorPost, visitorPre, context) {          }*/             return ret;             }                 }                     ret = ret.concat(ast[i]);                 else {                 }                             // }                             // }                             ret = ret.concat(createNewStatement( ast[i].expression ));                         //   if (node.left.property.name === "innerHTML") {                     //if (node.type == "AssignmentExpression" ) {                     ret = ret.concat(ast[i]);                 if ( ( ast[i].type == "ExpressionStatement") ) {             for (var i=0; i<ast.length; i++) {             var ret=[];         function instrumentUnary(node, ast) { ad     �     S       {  :    �  |  T  	  �  �  :  �  �  �  F     �  �  \    �
  �
  Q
  
  
  �	  ~	  X	  -	  �  �  [  A  +    �  �  �  x  X  <  .  -  �  �  �  �  f  =    �  �  �  m  [    �  �  �  t  a  `  _  %    �  �  {  U  ?      
  �  �  �  ^  8  "      �  �  �  �                                                     while (s !== null) {                     var s = this;                 Scope.prototype.addArguments = function() {                  };                     }                         s = s.parent;                         s.hasEval = true;                     while (s !== null) {                     var s = this;                 Scope.prototype.addEval = function() {                  };                     return null;                     }                         s = s.parent;                             return s.vars[name];                         if (HOP(s.vars,name))                     while (s !== null) {                     var s = this;                 Scope.prototype.hasVar = function(name) {                   };                     }                         //this.funLocs[name] = loc;                     if (type === 'defun') {                     this.vars[name] = type;                 Scope.prototype.addVar = function(name, type, loc) {                 }                     this.parent = parent;                     this.hasArguments = false;                     this.hasEval = false;                     //this.funLocs = {};                     this.vars = {};                 function Scope(parent) {             function addScopes(ast) {              */             http://tobyho.com/2013/12/02/fun-with-esprima/             /* The following  tutorial is good for understanding the scope variables               }                 return ret;                     ret = node;                 else                 }                     ret = visitorPost[type](node, context);                 if (visitorPost && HOP(visitorPost, type) ) {                 }                     }                         }                                     node[key] = transformAst(child, visitorPost, visitorPre, newContext);                                     }                                         newContext = CONTEXT.RHS;                                     else {                                     }                                         newContext = CONTEXT.IGNORE;                                     else if (context === CONTEXT.INC) {                                          newContext = CONTEXT.IGNORE;                                     else if (context===CONTEXT.OEXP3)                                     }                                         newContext = CONTEXT.OEXP3;                                     else if (context===CONTEXT.OEXP2 && key === 'value') {                                     }                                         newContext = CONTEXT.IGNORE;                                     else if (context===CONTEXT.OEXP2 && key === 'key') {                                     }                                         newContext = CONTEXT.OEXP2;                                     else if (context===CONTEXT.OEXP) {                                     }                                         newContext = CONTEXT.OEXP;                                     else if (type === 'ObjectExpression' && key === 'properties') {                                     }                                         newContext = CONTEXT.IGNORE;                                     else if (context === CONTEXT.PARAMS) {                                     }*/                                     CONTEXT.INC;                                 /*           else if (type === 'UpdateExpression' && key === 'argument') {                                 }                                     newContext = CONTEXT.PARAMS;                                 else if ( ((type === 'FunctionExpression' || type === 'FunctionDeclaration') && key === 'params') ){ ad     �     \       �  �  �  �  �  I         �  �  �  �  �  c  b  7    �  �  \    �  �  x  3    �  �  e  !    �
  �
  �
  �
  t
  b
  a
  4
  �	  �	  �	  �	  |	  [	  I	  H	  	  �  �  �  p  :  �  �  v  ;      �  �  v  7      �  �  �  �  Q  0    �  �  �  =  <  �  �  �  �  �  p  G    �  �  ?  -  �  �  �                                                   indent: { adjustMultilineComment: true}                   var codegenerateoptions = { comment: true, format: {                  }                     ast = transformAst(ast, visitorRRPost, visitorRRPre,  CONTEXT.RHS);                     addScopes(ast);                     //asttemp = transformAst(asttemp, visitorRRPost, visitorRRPre,  CONTEXT.RHS);                     //addScopes(asttemp);                     //var asttemp = ast;                 if (this.options.PARSING_MODE === "PARSE") {                   ast = escodegen.attachComments(ast, ast.comments, ast.tokens);                  var ast = esprima.parse(code, parseoptions);                  var parseoptions = { comment: true, range: true, tokens: true };                    //                  tokens: true, raw: true};                 //var parseoptions = { comment: true, loc: true, range: true,                  }                     return code;                 if (this.options.PARSING_MODE === "MINIFIED" ) {             this.instrument = function(code) {              }                             transformAst(ast, visitorPost, visitorPre);                              }                                 'FunctionExpression': popScope                                 'FunctionDeclaration': popScope,                                 'Program': popScope,                             var visitorPost = {                              }                                 'CatchClause': handleCatch                                 'VariableDeclarator': handleVar,                                 'FunctionExpression': handleFun,                                 'FunctionDeclaration': handleFun,                                 'Program': handleFun,                 var visitorPre = {                  // case where a variable is declared globally                 // 'AssignmentExpression' if we want to handle the                 //In the following, we should add:                  }                     return node;                     currentScope = currentScope.parent;                 function popScope(node) {                  }                     currentScope.addVar(node.param.name, "catch");                 function handleCatch(node) {                  }                     currentScope.addVar(node.id.name, "var");                 function handleVar(node) {                  }                     }                         })                             currentScope.addVar(param.name, "arg");                         MAP(node.params, function(param) {                         }                             currentScope.addVar(node.id.name, "lambda");                         if (node.id !== null) {                     } else if (node.type === 'FunctionExpression') {                         })                             currentScope.addVar(param.name, "arg");                         MAP(node.params, function(param) {                         oldScope.addVar(node.id.name, "defun", node.loc);                     if (node.type === 'FunctionDeclaration') {                     node.scope = currentScope;                     currentScope = new Scope(currentScope);                     var oldScope = currentScope;                 function handleFun(node) {                  var currentScope = null;                   };                     return this.hasArguments;                 Scope.prototype.usesArguments = function() {                  };                     return this.hasEval;                 Scope.prototype.usesEval = function() {                  };                     }                         s = s.parent;                         s.hasArguments = true; ad  �  �     6       �  �  `  L    �  �  �  c  @  -      �  �  N  (      �  �  �  �  �  =      �  �  _  �
  �
  �
  �
  y
  X
  �	  �	  �	  �	  o	  $	  �  �  g  $    �  �  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            function getPrope    function getPropertyAsAst(ast) {       }         }                 return node;              }                 node.right = ret;                 ret = instrumentAccumulationPoint(node, ReUseLId);                 // right one.                 // left side and the object on the right side by wrapping the                  // TODO in script to process data: connect the container on the                 // get the iid of the left side and use that for the right             if ( (thatModule.options.ACCUMULATION_POINT==1) && (rightType===true)) {              }                 node.left = ret;                 ret = wrapGetPutField(node.left, logFunctionName(loggerLib.consts.logPutFieldDot));                 ReUseLId = true;             else if (thatModule.options.WRITE_INST===1) {             }                 }                     node.left = ret;                     ret = wrapGetPutField(node.left, logFunctionName(loggerLib.consts.logPutDotNull));                 if (thatModule.options.RECORD_RIGHT_NULL===1) {                 rightType = false;             if ((node.right.type==="Literal")&&(node.right.value===null))  {                          // it is set to Null             //TODO: remove the following, later add support for the case that             var rightType=true;             var ReUseLId = false;          } else {  //a.b =              return node;                  }                  }                     node.right = ret;                     ret = instrumentIdentifierSetNull(node);                     if ((node.right.type==="Literal")&&(node.right.value===null))  {              if (thatModule.options.RECORD_RIGHT_NULL===1) {               }                  }                  node.right = ret;                  ret = instrumentWriteToIdentifier(node);                 else {                 }                 if ((node.right.type==="Literal")&&(node.right.value===null)) {              if (thatModule.options.WRITE_INST===1) {             // }                //    node.right = ret;             //    ret = instrumentGlobalVariableReference(node);             //if (thatModule.options.GLOBAL_VAR_REF===1) { 