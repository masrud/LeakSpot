b0VIM 7.3      ��JT�B� �F  masoomeh                                masoomeh-ThinkPad                       ~masoomeh/Research/DevelopedTools/HttpsProxy/lib/profilerLib.js                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              utf-8 3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp	           C                     	       $       E                     6       f              
              �                     8       �                     1       �                     h                           d       �                    "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad  �  �     C       �  �  �  �  w  \  7      �  v  d  F  E  /  
  �  �  �  �  l  H  $    �  �  �  �  q  Q  -  
  �  �  �  |  Z  @    �
  �
  �
  �
  �
  �
  l
  <
  
  �	  �	  �	  N	  -	  	  �  R  4  �  �  �    [  J  ?    �  �  �  �  p  :    �  �  �  y  I  7  
  �  �  d  @  2  (  �  �  �  y  Q  ,    �  �  �  w  8      �  �  �                  return function() {         function wrapFunc(func, type) {         }             }                 return returnvalue;                 var returnvalue = func.apply(this, arguments);                 arguments[0] = xhr.responseText;                 }                     console.log(xhr.responseText);                     console.log("response");                 {                 if (xhr.status==200)                 xhr.send(arguments[0]);                 xhr.open("POST", "/HTMLData", false);                 var xhr = new XMLHttpRequest();             return function() {         function wrapWrite(func, type) {         }             }                 return returnvalue;                 var returnvalue = func.apply(this, arguments);                 arguments[0] = xhr.responseText;                   //console.log(typeof arguments[0]);                 //console.log(arguments[0]);                 }                     //TODO: update arguments[0]                     //console.log(xhr.responseText);                     console.log("response");                 {                 if (xhr.status==200)                 xhr.send(arguments[0]);                 xhr.open("POST", "/HTMLData", false);                 var xhr = new XMLHttpRequest();                 //console.log(arguments);                             if (evalMonitor===1) {             return function() {         function wrapEval(func) {         }              }                    return returnvalue;                 }                     }                         logLine(line);                             line = [constants.UNKNOWN, type, res1.oid, findproto(this),"\n"].join();                          else                              line = [constants.UNKNOWN, type, res1.oid, findproto(this), res2.oid, findproto(arguments[0]), "\n"].join();                          if (res2.stat>0)                      if (res1.stat>0) {                     var line="";                     var res2 = addObjectId(arguments[0]);                     var res1 = addObjectId(this);                 if (Logging === 1) {                 var returnvalue=func.apply(this, arguments);             return function() {         function wrapArrayPushPop(func, type) {     if (typeof window !=='undefined') {     this.consts = constants;      };         UNKNOWN : "-1"         logWriteUndefinedNull : "LWUNull",         logWriteUndefined : "LWU",          logWriteNull : "LWNull",         logWrite : "LWR",         logReadUndefined : "LRU",         logRead : "LRE",         logRightSidePutDot : "LRSP",         logRightSidePutBracket : "LRPE",         logPutBracketNull : "LPENull",         logPutDotNull : "LPDNull",         logPutFieldBracket : "LPE",         logPutFieldDot : "LPD",         logMethodCall : "LMC",         logLiteral : "T",         logNewFunction : "LNF",         logNewObject : "LNE",         logUndefined : "I",         logGetFieldDot : "LGD",         logGetFieldBracket : "LGE",         logFuncDeclaration : "LFD",         logFuncCall : "LFC",         logArrayPop: "ArrPop",         logArrayPush: "ArrPush",         objectCreate : "objCr",         WrapWrite : "WrapWrite",         DOMCreateElement : "CRElem",     var constants = {      var INTERVALTIME = 60000;     this.TMPS={};      var MAX_BUF_SIZE = 23107200;  //131072   1024*64 = 65635     var ReferenceCreation = 1 //This should be 1 if want to measure just beautify     var DOMLogging = 1;     var evalMonitor = 0;     var Logging = 1; //On==1, Off==0     var COMMUNICATION = 1;     var objectId = 1; JSProf = new ( function() {  //eval, document.write.... //TODO: We have used function wrapping to cover the cases: ad  �
  �     "       �  �  d  Z  D  >  =  �  �  �  �    �  �  �  �  �  �  {  `  7    �  �  �  s  i  S  M    �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          })();     }         return right;         //This never generate anythings, since left is undefined and right is null     this[this.consts.logWriteUndefinedNull] = function (iid, left, right) {     }         return right;         }             }                 logLine(line);                 line = [iid, constants.logWriteNull, res.oid, findproto(left), "\n"].join();             if (res.stat > 0 ) {             var line="";             var res = addObjectId(left);         if (Logging===1) {     this[ this.consts.logWriteNull ] = function (iid, left, right) {       }         return right;         }             }                 logLine(line);                    var line = [iid, constants.logWriteUndefined, resRight.oid,findproto(right), "\n"].join();             if ( resRight.stat > 0 ) {             var resRight = addObjectId(right);         if (Logging===1) {     this[ this.consts.logWriteUndefined ] = function(iid, left, right) {      }         return right;         }              logLine(line);                                line = [iid, constants.logWrite, constants.UNKNOWN , resleft.oid, findproto(left), "\n"].join(); ad  �  �     1       �  s  r  R    �  �  �  �  W  7  �  �  s  \  �  �  �  �  w  e  :  9  $  �  �  �  �  �  �  b  \  "  �
  �
  �
  �
  z
  
  �	  �	  �	  �	  �	  ;	  	  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        eval = wrapEval(eval);             var prop = eval("baseobj."+propname);             eval = originalEval;         if ( Logging === 1 ) {     this[ this.consts.logGetFieldDot ] = function(iid, baseobj, propname) {     }         }            logLine(line);                line = [iid, action, res1.oid, findproto(base), "\n"].join();              else                  line = [iid, action, res1.oid, findproto(base), res2.oid, findproto(prop), "\n"].join();             if (res2.stat > 0 )              var res2 = addObjectId(prop);             var line="";         if ( res1.stat > 0) {         var res1 = addObjectId(base);     function generateGetPutLog(iid, action, base, prop) {     }                 sendToServer(line, false);                if (line.length > 0)         if (COMMUNICATION===1)     function logLine(line) {     }         }             return {stat:-1, oid: -1};         } catch(e) {                  return {stat:-1, oid: -1};             else              }                 }                     return {stat:1, oid: oidval};                     //var oidval = obj.__objectID__ ;                     var oidval = Object.getOwnPropertyDescriptor(obj, "__objectID__").value;                 else {                 }                     return {stat: 2 , oid:objidvalue};                     Object.defineProperty(obj, "__objectID__", { enumerable: false, value: objidvalue, writable: false });                     objectId++;                     var objidvalue = objectId + "" +  SUFFIX;                     }                             SUFFIX = suffix;                     else {                          SUFFIX = 'S2';                     if (typeof window === 'undefined')                     var SUFFIX;                      //if sizing information is required.                     //TODO: If enumerable is false, can it be seen by heap snapshot ad  u  q     8       �  �  �  m  '    �  �  �  �  M  *    �  �  �  �  �  G      �  �  e  ,            �  �  �  �    �
  �
  �
  �
  a
  `
  =
  +
  
  �	  �	  �	  �	  �	  �	  �	  }	  2	  �  �  q  [  Z  :    �  �  �  }  ?    �  m  [  D  �  �  �  �  �  X  W  B        �  �  �  �  z  @    �  �  �  �  /    �  �  �  �  Y  :    �  �                              eval = wrapEval(eval);             var prop = eval("baseobj."+propname);             eval = originalEval;         if ( Logging === 1 ) {     this[ this.consts.logGetFieldDot ] = function(iid, baseobj, propname) {     }         }            logLine(line);                line = [iid, action, res1.oid, findproto(base), "\n"].join();              else                  line = [iid, action, res1.oid, findproto(base), res2.oid, findproto(prop), "\n"].join();             if (res2.stat > 0 )              var res2 = addObjectId(prop);             var line="";         if ( res1.stat > 0) {         var res1 = addObjectId(base);     function generateGetPutLog(iid, action, base, prop) {     }                 sendToServer(line, false);                if (line.length > 0)         if (COMMUNICATION===1)     function logLine(line) {     }         }             return {stat:-1, oid: -1};         } catch(e) {                  return {stat:-1, oid: -1};             else              }                 }                     return {stat:1, oid: oidval};                     var oidval = Object.getOwnPropertyDescriptor(obj, "__objectID__").value;                 else {                 }                     return {stat: 2 , oid:objidvalue};                     Object.defineProperty(obj, "__objectID__", { enumerable: false, value: objidvalue, writable: false });                     objectId++;                     var objidvalue = objectId + "" +  SUFFIX;                     }                             SUFFIX = suffix;                     else {                          SUFFIX = 'S2';                     if (typeof window === 'undefined')                     var SUFFIX;                                        if (!Object.prototype.hasOwnProperty.call(obj, "__objectID__")) {                 //if ( obj.__objectID__ === undefined  ) {             (obj !== null)&&(obj !== undefined)) {              if (((typeof obj === 'object')||(typeof obj === 'function'))&&         try {     function addObjectId (obj) {     }         }             return "";         } catch(e) {             return "";             }                 return tname;                 }                     tname += name;                          name = "0";                     if (name=="")                     var name = objprototype.constructor.name;                  if (objprototype!==null) {                 var objprototype =  Object.getPrototypeOf(obj); // Catch since sometime these are from two origins TODO             if ( (obj!== null) || (obj !== undefined) ) {         try{         var tname="";     function findproto(obj) {      }         },false);              }                 logLine("\nemptybuffer--"+suffix+"\n" );                 //sendToServer("\nemptybuffer--"+suffix+"\n", true);             if (event.data.type && (event.data.type == "FROM_CONTENT")) {             }                    return;             if (event.source != window) {         window.addEventListener('message',function(event) {         }              }                 inbrowserbufferSize = 0;                 console.log("errror ...........sending data");                 inbrowserbuffer = "";                 intervalOn = true;                 //console.log("error transfering "+ xhrBUFFER.status);             else {             }                 inbrowserbufferSize = 0;                 inbrowserbuffer = "";                 intervalOn = true;             if (xhrBUFFER.status == 200 || xhrBUFFER.status == 304) {             xhrBUFFER.send(inbrowserbuffer);             xhrBUFFER.open("POST", "/POST_MONITORING_DATA", false);             }*/                 } ad     �     h       �  �  �  �  �  5    �  �  �  �  S  6  
  �  �  q  c  Y  (  �  �  S  B  6  0  /  �  �  �  �  0    �
  �
  �
  �
  �
  �
  p
  B
  �	  �	  �	  �	  r	  <	  	  �  �  �  �  |  v  u    �  �  �  �  �  B  %    �  �  �  x  _  Q    �  �  �  �  �  d    �  �  �  �  �  s  R  �  �  �  �  �  �  m  S    �  �  �  �  K  7  1  0  �  �  �                             if (Logging===1) {     this[ this.consts.logNewObject ] = function(iid, obj, objtype ) {      }         return obj;            generateRightSide(iid, constants.logRightSidePutDot, obj);         if (Logging===1)      this[ this.consts.logRightSidePutDot ]  = function(iid, obj) {     }         return obj;             generateRightSide(iid, constants.logRightSidePutBracket, obj);         if (Logging===1)      this[ this.consts.logRightSidePutBracket ] = function(iid, obj) {      }         }             }                 logLine(line);                     var line = [iid, action, res.oid, findproto(baseobj), res.oid, "\n"].join();             if (res.stat > 0 ) {             var res = addObjectId(baseobj);         if (Logging===1) {     function generateRightSide(iid, action, baseobj ) {      }         return baseobj;             generateGetPutLog(iid, constants.logPutBracketNull, baseobj, realobj);         if (Logging === 1)      this[ this.consts.logPutBracketNull ] = function(iid, baseobj, propname, realobj ) {      }         return baseobj;         }             generateGetPutLog(iid, constants.logPutDotNull, baseobj, realobj);             }             } catch(e) {                 eval = wrapEval(eval);                 realobj = eval("baseobj."+propname);                  eval = originalEval;             try {             var realobj;         if (Logging === 1) {     this[ this.consts.logPutDotNull ] = function(iid, baseobj, propname) {      }         return baseobj;            generateGetPutLog(iid, constants.logPutFieldBracket, baseobj, realobj);         if (Logging === 1)      this[ this.consts.logPutFieldBracket ] = function(iid, baseobj, propname, realobj ) {      }         return baseobj;         }             generateGetPutLog(iid, constants.logPutFieldDot, baseobj, realobj);             }             } catch(e) {                 eval = wrapEval(eval);                 realobj = eval("baseobj."+propname);                  eval = originalEval;             try {             var realobj;              //that this is an add of property.             //check to see if obj[name] already exist or not! if not this means             //To distinguish add from update:         if (Logging === 1) {     this[ this.consts.logPutFieldDot ] = function(iid, baseobj, propname) {      }         return func;         }             }                 logLine(line);                     var line = [iid, constants.logFuncCall, res.oid, "\n"].join();              if (res.stat>0) {             var res = addObjectId(func);         if (Logging === 1) {     this[ this.consts.logFuncCall ] = function(iid, func, isConstructor) {      }         }*/             }                    line += iid+ " Dec " + res2.oid + " +prototype" + " " + "\n";              if (res2.stat > 0){             var res2 = addObjectId(funcobj.prototype); //This is not needed for memory leak detection         /*if ( funcbj.prototype != undefined ) {         }             }                 logLine(line);                      var line = [iid,constants.logFuncDeclaration,res.oid,"\n"].join();              if ( res.stat > 0) {             var res = addObjectId(funcobj);         if (Logging === 1) {     this[ this.consts.logFuncDeclaration ]  = function (iid, funcobj, isCtr) {          }         return baseobj;             generateGetPutLog(iid, constants.logGetFieldBracket, baseobj, realobj);         if (Logging === 1)      this[ this.consts.logGetFieldBracket ] = function(iid, baseobj, prop, realobj) {      }         return baseobj;         }             generateGetPutLog(iid, constants.logGetFieldDot, baseobj, prop); ad  >   �     d       �  �  �  �    �  �  j  \  R  >  8  7  �  �  �  �  ;        �  �  �  �  �  x  "  �  �  �  �  �  `  R  ?    �
  �
  �
  �
  �
  k
  3
  	
  �	  R	  @	  *	  �  �  �  ~  f  `  _           �  �  �  �  r  W  /    �  �  p  Z    �  �  �  �  �  �  m  R  *    �  �  t  j  V  P  O    �  �  �  {  9  �  �    �  �                                                                             else if ( ( resleft.stat > 0 ) )                   line = [iid, constants.logWrite, resright.oid, findproto(right), constants.UNKNOWN, "\n"].join();              else if ( (resright.stat > 0 ) )                   line = [iid, constants.logWrite, resright.oid, findproto(right), resleft.oid, findproto(left), "\n"].join();              if ( (resright.stat > 0 ) && ( resleft.stat > 0 ) )               var resright = addObjectId(right);              var resleft = addObjectId(left);              var line="";         if (Logging===1) {     this[ this.consts.logWrite ] = function (iid, left, right) {      }         return obj;         }             }                 logLine(line);                    var line = [iid, constants.logReadUndefined, res.oid, findproto(obj), "\n"].join();             if ( res.stat > 0 ) {             var res = addObjectId(obj);         if (Logging===1) {     this[ this.consts.logReadUndefined ] = function (iid, obj) {       }         return obj;         }             }                 logLine(line);                     line = [iid,constants.logRead,res.oid, findproto(obj), "\n"].join();                 else                      line = [iid,constants.logRead,res.oid, findproto(obj), "NEW","\n"].join();                  if (res.stat === 2)              var line="";             if (res.stat > 0 ) {             var res = addObjectId(obj);         if (Logging===1) {     this[ this.consts.logRead ] = function(iid, obj) {      }             return val;      this[ this.consts.logUndefined ] = function (val) {          }         return obj;     this[this.consts.logLiteral] = function (iid, obj, type) {      }         return baseobj;         }              }                 logLine(line);                     line = [iid,constants.logMethodCall, resBase.oid,findproto(baseobj), methodname, "\n"].join();                  else                  }                             resMethod.oid, findproto(methodobj), methodname, "\n"].join();                      line = [iid,constants.logMethodCall, resBase.oid, findproto(baseobj),                  if (resMethod.stat > 0) {                 var resMethod = addObjectId(methodobj);             var line="";             if (resBase.stat>0) {             var resBase=addObjectId(baseobj);             eval = wrapEval(eval);              }                 methodobj = eval("baseobj."+methodname);             else {             }                 methodobj = eval("baseobj[methodname]");             if (type !== undefined) {             eval = originalEval;              var methodobj;             // push/pop or call/apply             // The methodname is used for finding the location in the code in case of         if (Logging===1) {      this[ this.consts.logMethodCall ] = function(iid, baseobj, methodname, type) {        }         return obj;         }             }                 logLine(line);                 var line = [iid, constants.logNewFunction, res.oid, "\n"].join();              if (res.stat>0) {             var res = addObjectId(obj);         if (Logging===1) {     this[ this.consts.logNewFunction ] = function(iid, obj, objtype ) {      }         return obj;         }             }                 logLine(line);                     line = [iid, constants.logNewObject, res.oid, objtype, findproto(obj), "\n"].join();                  else                             line = [iid, constants.logNewObject, res.oid, objtype, findproto(obj), "SURPRISE\n"].join();                 if (res==1)                 var line="";             if (res.stat>0) {             var res = addObjectId(obj); ad    	     6       �  �  u  O  �  �  �  �  �  o  b    �  �  '      �  �  G  &    �  p  o  :    �
  K
  
  �	  Y	  6	  5	  �  �  {  A  �  �  �  �  �  �  f  D       �  �  �  7    	  �  �  �  W  -    �  �  �  �  �  <  �  �  �  �  y  9    �  �  N  #    �  �  z  d                          }                         intervalOn = true;                         console.log("error transfering "+ xhrBUFFER.status);                     else {                     }                         intervalOn = true;                     if (xhrBUFFER.status == 200 || xhrBUFFER.status == 304) {                 if (xhrBUFFER.readyState == 4) {             /*xhrBUFFER.onreadystatechange = function() {             var xhrBUFFER = new XMLHttpRequest();             //async: true (asynchronous) or false (synchronous)             intervalOn = false;         function sendInterval() {          // is not set to true when it is needed.          // not being executed at the time I'm expecting. Therefore intercalOn         // because onreadystatechange is a callback function, it is         }             window.setInterval(sendToServerPeriodically, INTERVALTIME);         if (COMMUNICATION === 1) {         }             }                 sendInterval();                 //console.log("*******");             if ( intervalOn &&  (inbrowserbufferSize > 0) ) {             //console.log("............."+intervalOn);         function sendToServerPeriodicall            //}                  }                 sendInterval();             if ( (inbrowserbufferSize >= MAX_BUF_SIZE) && (intervalOn) ) {             inbrowserbufferSize += msg.length;             inbrowserbuffer += msg;         function sendToServer(msg, imm ) {         var intervalOn = true;         var inbrowserbufferSize = 0;         var inbrowserbuffer = "";     if (typeof window !== 'undefined') {     }             }, 2000); } );                  logLine(line);                      xhr.send("load time = "+ loadtime +" location origin : " + window.location.origin + "\n" );                     xhr.open("POST", "/LOADDATA", false);                     var xhr = new XMLHttpRequest();                 //It does not add it to the buffer                 //Send the load time of a page instantly to the proxy to be logged                  console.log(line);                 var line = "load time = "+ loadtime +" location origin : " + window.location.origin + "\n";                 console.log("load time in seconds" + loadtime);                 //Therefore, we are diving by 1000 to have in seconds                 //Time returned by window.performance.timing is in milliseconds.                 var loadtime = (window.performance.timing.loadEventEnd - window.performance.timing.navigationStart)/1000;             setTimeout(function() {         window.addEventListener('load', function() {          Document.prototype.createElement = wrapFunc(Document.prototype.createElement, constants.DOMCreateElement);             eval = wrapEval(eval);         if (evalMonitor === 1 )         var originalEval = eval;         //HTMLDocument.prototype.write = wrapWrite( HTMLDocument.prototype.write, constants.WrapWrite);           //add Call Apply, since the first argument of this function is access to an object.         //TODO:         }             //Array.prototype.pop  = wrapArrayPushPop( Array.prototype.pop, constants.logArrayPop );             Array.prototype.push = wrapArrayPushPop( Array.prototype.push, constants.logArrayPush );         if ( ReferenceCreation == 1 ) {         Object.create = wrapFunc(Object.create, constants.objectCreate);         }                }                    return ret;                 }                     }                         logLine(line);                         var line = [constants.UNKNOWN, type,res.oid, findproto(ret), "\n"].join();                      if (res.stat>0) {                     var res = addObjectId(ret);                 if (DOMLogging===1) {                 var ret=func.apply(this, arguments); ad  �	  {
     $       �  �  u  ;    �  �  �  f  2    �  �  |  j  +    �  �  �  �  v  @    �  �  �  �  o  >  �
  �
  �
  �
  �
  {
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 return function() {         function wrapFunc(func, type) {         }             }                 return returnvalue;                 var returnvalue = func.apply(this, arguments);                 arguments[0] = xhr.responseText;                 }                     console.log(xhr.responseText);                     console.log("response");                 {                 if (xhr.status==200)                 xhr.send(arguments[0]);                 xhr.open("POST", "/HTMLData", false);                 var xhr = new XMLHttpRequest();             return function() {         function wrapWrite(func, type) {         }             }                 return returnvalue;                 var returnvalue = func.apply(this, arguments);                 }                     arguments[0] = xhr.responseText;                       //console.log(typeof arguments[0]);                     //console.log(arguments[0]);                     }                         //TODO: update arguments[0]                         //console.log(xhr.responseText);                         console.log("response");                     {                     if (xhr.status==200)                     xhr.send(arguments[0]);                     xhr.open("POST", "/HTMLData", false);                     var xhr = new XMLHttpRequest();                     //console.log(arguments);                     //console.log(this); ad  �
  `            �  �  �  S  )  	  �  �  �  �  |  8  �  �  �  �  u  5    �  �  J    	  �  �  v  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                         intervalOn = true;                         console.log("error transfering "+ xhrBUFFER.status);                     else {                     }                         intervalOn = true;                     if (xhrBUFFER.status == 200 || xhrBUFFER.status == 304) {                 if (xhrBUFFER.readyState == 4) {             /*xhrBUFFER.onreadystatechange = function() {             var xhrBUFFER = new XMLHttpRequest();             //async: true (asynchronous) or false (synchronous)             intervalOn = false;         function sendInterval() {          // is not set to true when it is needed.          // not being executed at the time I'm expecting. Therefore intercalOn         // because onreadystatechange is a callback function, it is         }             window.setInterval(sendToServerPeriodically, INTERVALTIME);         if (COMMUNICATION === 1) {         }             }                 sendInterval();                 //console.log("*******");             if ( intervalOn &&  (inbrowserbufferSize > 0) ) {             //console.log("............."+intervalOn);         function sendToServerPeriodically() {         } 